

o intro
        - vip core, supports 3 version of axi(3,4,lite)
        - unencrypted SV source[synthesizeable RTL?] ( difference b/w IP & VIP ?)
        - m_axi, s_axi & pass-thru which acts as monitor. ( by using this VIP, we are generating transactions ?)

o

